`timescale 1ns/1ns

module alu();

endmodule

module ramS();

endmodule

module instructionRam();

endmodule

module registerBank();

endmodule

module vCoreZero();

endmodule